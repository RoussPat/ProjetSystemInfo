`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:53:14 04/19/2020 
// Design Name: 
// Module Name:    registre 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module registre(
    input [3:0] A,
    input [3:0] B,
    input [3:0] W,
    input Write,
    input [7:0] DATA,
    input RST,
    input CLK,
    output [7:0] QA,
    output [7:0] QB
    );


endmodule
